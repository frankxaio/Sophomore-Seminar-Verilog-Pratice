`timescale 1ns / 1ps

module test_bench;
	
	reg [9499:0] A;
	reg [18999:0] B;
	
	wire [3799:0] Answer;
	
	Calculator calculator(.A(A), .B(B), .Result(Answer));
	
	initial begin
		
		//Initial inputs
		A={-19'd188, 19'd168, 19'd95, -19'd141,
			 19'd50, -19'd182, -19'd216, 19'd26, -19'd185, 19'd64, 19'd85, -19'd8, 19'd201, 19'd192, -19'd3, 19'd247, 19'd129, 19'd244, 19'd67, -19'd45, 19'd23, 19'd70, 19'd32, -19'd61, 19'd214, -19'd207, 19'd133, 19'd249, -19'd67, -19'd144, -19'd7, 19'd87, -19'd79, 19'd67, -19'd197, 19'd69, -19'd177, -19'd55, 19'd166, 19'd146, 19'd72, -19'd137, 19'd252, -19'd168, 19'd185, 19'd148, 19'd160, -19'd57, 19'd170, 19'd195, 19'd182, -19'd193, -19'd32, -19'd45, 19'd189, -19'd153, 19'd210, 19'd176, -19'd5, -19'd113, 19'd245, 19'd77, -19'd163, -19'd69, 19'd76, 19'd187, -19'd126, 19'd234, -19'd127, -19'd208, -19'd114, -19'd244, 19'd101, 19'd53, 19'd91, -19'd247, -19'd59, 19'd220, 19'd218, 19'd231, 19'd185, -19'd26, -19'd63, 19'd110, 19'd221, 19'd93, -19'd215, -19'd29, 19'd153, -19'd151, -19'd45, -19'd158, 19'd9, -19'd238, -19'd40, -19'd69, -19'd42, 19'd63, -19'd31, -19'd187, -19'd26, -19'd88, 19'd159, -19'd9, 19'd33, 19'd248, -19'd45, 19'd233, 19'd137, 19'd15, 19'd41, -19'd46, 19'd249, -19'd203, -19'd119, 19'd231, -19'd185, 19'd84, 19'd42, -19'd193, -19'd10, 19'd145, 19'd173, -19'd66, 19'd141, -19'd135, -19'd9, 19'd62, 19'd240, -19'd137, -19'd98, 19'd95, 19'd137, 19'd172, 19'd91, 19'd134, -19'd197, 19'd101, 19'd84, 19'd248, -19'd245, 19'd170, 19'd74, 19'd114, -19'd152, -19'd37, -19'd10, -19'd46, 19'd156, -19'd79, 19'd226, -19'd125, 19'd193, -19'd253, 19'd52, -19'd224, -19'd206, -19'd50, -19'd140, -19'd65, -19'd229, 19'd252, -19'd62, 19'd104, -19'd170, -19'd206, 19'd244, 19'd251, 19'd194, -19'd103, 19'd116, 19'd217, 19'd69, -19'd252, 19'd231, -19'd109, 19'd204, 19'd41, 19'd228, -19'd80, -19'd204, -19'd160, -19'd18, -19'd20, 19'd72, -19'd140, 19'd210, -19'd124, 19'd196, -19'd200, 19'd214, 19'd178, -19'd221, -19'd237, -19'd31, -19'd157, -19'd152, -19'd114, -19'd244, -19'd217, -19'd172 ,19'd53 ,-19'd173 ,19'd203 ,-19'd129 ,19'd120 ,19'd194 ,-19'd229 ,19'd65 ,19'd32 ,-19'd16 ,-19'd242 ,19'd93 ,-19'd146 ,19'd132 ,-19'd61 ,19'd228 ,-19'd75 ,-19'd34 ,-19'd82 ,-19'd150 ,-19'd21 ,-19'd208 ,19'd252 ,19'd224 ,-19'd87 ,19'd43 ,19'd221 ,-19'd170 ,19'd40 ,-19'd39 ,-19'd67 ,19'd185 ,19'd116 ,-19'd121 ,-19'd91 ,19'd178 ,-19'd87 ,19'd33 ,-19'd25 ,19'd191 ,-19'd88 ,19'd122 ,19'd189 ,19'd88 ,-19'd141 ,19'd151 ,-19'd102 ,19'd34 ,-19'd74,-19'd234 ,-19'd106 ,-19'd9 ,19'd93 ,19'd213 ,19'd197 ,19'd204 ,-19'd168 ,19'd130 ,19'd17 ,19'd186 ,19'd116 ,19'd128 ,-19'd36 ,-19'd40 ,-19'd243 ,19'd242 ,-19'd136 ,-19'd49 ,-19'd195 ,19'd71 ,19'd106 ,19'd251 ,19'd200 ,19'd215 ,-19'd129 ,-19'd57 ,19'd60 ,-19'd179 ,19'd6 ,19'd81 ,19'd229 ,19'd89 ,-19'd90 ,-19'd32 ,19'd193 ,19'd195 ,19'd153 ,19'd85 ,19'd22 ,19'd203 ,-19'd89 ,-19'd45 ,-19'd168 ,19'd252 ,-19'd116 ,19'd10 ,-19'd230 ,-19'd62 ,-19'd55,19'd230 ,19'd229 ,-19'd90 ,-19'd104 ,19'd216 ,19'd184 ,19'd56 ,-19'd73 ,19'd206 ,-19'd86 ,-19'd205 ,-19'd187 ,-19'd233 ,19'd24 ,19'd236 ,-19'd14 ,19'd181 ,19'd146 ,-19'd85 ,19'd238 ,-19'd147 ,19'd199 ,-19'd166 ,19'd58 ,-19'd220 ,19'd173 ,-19'd203 ,19'd107 ,-19'd34 ,19'd61 ,19'd168 ,-19'd195 ,19'd84 ,19'd216 ,19'd88 ,-19'd75 ,-19'd243 ,19'd166 ,-19'd48 ,19'd86 ,-19'd192 ,-19'd37 ,19'd5 ,-19'd50 ,19'd184 ,-19'd162 ,-19'd39 ,-19'd203 ,19'd92 ,-19'd192,-19'd144 ,-19'd251 ,19'd228 ,-19'd126 ,-19'd12 ,19'd199 ,-19'd249 ,-19'd124 ,19'd102 ,19'd243 ,19'd28 ,19'd59 ,19'd229 ,19'd2 ,19'd213 ,-19'd47 ,-19'd123 ,-19'd137 ,19'd195 ,19'd6 ,19'd72 ,-19'd114 ,-19'd230 ,-19'd164 ,-19'd169 ,-19'd89 ,-19'd34 ,19'd6 ,-19'd251 ,-19'd82 ,19'd232 ,-19'd64 ,19'd221 ,-19'd227 ,19'd95 ,19'd75 ,19'd30 ,19'd138 ,-19'd14 ,-19'd66 ,-19'd12 ,-19'd64 ,-19'd122 ,19'd87 ,-19'd98 ,19'd229 ,19'd120 ,19'd106 ,19'd103 ,-19'd232,-19'd101 ,-19'd148 ,-19'd98 ,19'd27 ,19'd70 ,-19'd213 ,19'd78 ,19'd247 ,19'd7 ,19'd165 ,-19'd217 ,19'd64 ,-19'd254 ,-19'd123 ,19'd92 ,19'd223 ,19'd49 ,-19'd7 ,-19'd136 ,-19'd227 ,-19'd105 ,19'd41 ,-19'd143 ,19'd131 ,19'd43 ,19'd84 ,19'd173 ,-19'd125 ,-19'd65 ,-19'd81 ,19'd112 ,19'd199 ,-19'd148 ,19'd173 ,19'd82 ,19'd63 ,19'd6 ,-19'd239 ,-19'd83 ,-19'd157 ,19'd39 ,-19'd56 ,-19'd189 ,-19'd106 ,19'd6 ,19'd228 ,-19'd69 ,19'd202 ,19'd68 ,19'd226,19'd116 ,19'd60 ,19'd55 ,19'd183 ,-19'd248 ,19'd201 ,-19'd208 ,-19'd55 ,-19'd159 ,-19'd225 ,19'd139 ,-19'd161 ,-19'd59 ,19'd46 ,19'd228 ,19'd148 ,-19'd3 ,19'd6 ,-19'd29 ,19'd106 ,-19'd11 ,19'd35 ,19'd222 ,-19'd75 ,-19'd113 ,-19'd70 ,-19'd240 ,-19'd251 ,19'd125 ,19'd15 ,19'd9 ,19'd99 ,-19'd49 ,19'd96 ,19'd249 ,19'd202 ,19'd162 ,19'd234 ,19'd192 ,19'd152 ,-19'd200 ,-19'd242 ,19'd211 ,19'd7 ,19'd148 ,19'd147 ,19'd48 ,-19'd136 ,19'd153 ,19'd200
		};
		B={-19'd43,19'd36,19'd26,-19'd9,
			19'd33,19'd19,-19'd2,-19'd33,-19'd7,19'd43,19'd0,19'd30,19'd49,-19'd47,19'd11,-19'd28,	19'd44,19'd32,-19'd13,19'd8,19'd17,19'd39,-19'd37,-19'd11,19'd45,19'd3,19'd39,19'd1,19'd12,-19'd22,-19'd5,-19'd26,19'd0,19'd17,19'd8,19'd21,19'd9,-19'd8,19'd38,19'd12,-19'd4,19'd42,-19'd24,-19'd11,-19'd38,19'd41,-19'd5,19'd47,-19'd50,19'd49,-19'd12,19'd7,-19'd7,-19'd20,-19'd23,19'd9,-19'd39,19'd15,-19'd36,-19'd9,-19'd47,19'd30,-19'd45,-19'd5,19'd2,19'd24,19'd21,19'd36,-19'd24,19'd26,19'd23,-19'd43,19'd36,-19'd15,19'd4,-19'd27,-19'd40,19'd15,-19'd23,19'd13,-19'd40,-19'd7,-19'd45,-19'd14,19'd3,-19'd42,-19'd17,19'd20,-19'd1,-19'd42,19'd23,19'd45,19'd42,-19'd39,19'd5,-19'd37,-19'd17,-19'd19,19'd14,-19'd33,19'd31,19'd49,19'd36,19'd1,19'd49,19'd3,-19'd11,-19'd5,-19'd40,19'd25,19'd1,19'd23,19'd28,-19'd12,-19'd8,19'd10,19'd39,-19'd4,19'd49,-19'd39,-19'd6,19'd21,-19'd8,19'd8,-19'd37,-19'd33,19'd22,-19'd29,-19'd31,-19'd4,19'd26,-19'd23,19'd11,-19'd15,-19'd45,-19'd33,19'd16,19'd28,19'd42,-19'd17,-19'd31,-19'd49,19'd40,19'd23,19'd21,19'd33,-19'd21,19'd25,-19'd34,-19'd25,-19'd35,-19'd34,19'd30,19'd29,-19'd21,19'd49,19'd36,-19'd32,19'd26,19'd10,-19'd10,-19'd15,-19'd46,-19'd36,-19'd29,19'd43,-19'd27,19'd27,-19'd28,-19'd16,-19'd19,-19'd13,-19'd5,-19'd41,19'd15,19'd23,-19'd28,-19'd20,19'd36,19'd37,-19'd13,19'd18,-19'd37,-19'd9,-19'd4,-19'd14,-19'd7,-19'd36,-19'd8,-19'd45,19'd8,19'd40,-19'd25,-19'd43,19'd46,-19'd34,19'd44,19'd2,-19'd33,19'd29,19'd32,-19'd3,19'd21,19'd32,19'd31,19'd44,-19'd38,-19'd10,-19'd42,-19'd23,19'd1,19'd8,-19'd12,-19'd34,19'd3,19'd0,-19'd14,19'd36,19'd26,19'd0,-19'd27,19'd14,19'd0,-19'd19,-19'd15,19'd15,19'd27,19'd19,19'd33,-19'd43,19'd29,19'd27,-19'd5,-19'd19,-19'd11,-19'd11,19'd1,19'd1,19'd10,19'd26,19'd18,19'd25,19'd18,19'd45,-19'd26,19'd30,-19'd44,-19'd38,-19'd1,19'd43,-19'd9,-19'd34,-19'd47,-19'd20,-19'd17,19'd7,19'd22,-19'd41,-19'd32,-19'd6,-19'd3,-19'd26,19'd1,19'd37,-19'd48,19'd49,19'd15,-19'd6,19'd0,-19'd18,19'd36,19'd16,-19'd34,19'd36,19'd0,19'd19,-19'd50,-19'd9,-19'd30,-19'd13,19'd9,19'd32,-19'd33,19'd31,19'd9,-19'd44,-19'd29,-19'd42,19'd37,19'd21,-19'd20,-19'd33,-19'd9,19'd12,-19'd49,19'd7,19'd50,19'd48,-19'd12,-19'd20,-19'd38,-19'd22,-19'd37,-19'd38,-19'd31,-19'd36,-19'd9,-19'd18,19'd11,-19'd48,19'd40,-19'd50,19'd16,19'd38,19'd28,-19'd18,19'd30,19'd24,-19'd2,19'd46,-19'd1,19'd2,19'd36,-19'd29,19'd21,19'd42,19'd24,-19'd24,19'd37,-19'd19,-19'd12,19'd49,-19'd28,19'd33,-19'd36,19'd22,19'd17,19'd32,-19'd21,-19'd44,19'd7,-19'd36,19'd41,19'd45,-19'd31,19'd46,19'd13,-19'd2,19'd4,-19'd44,19'd28,-19'd4,-19'd18,-19'd5,-19'd13,-19'd47,-19'd25,19'd46,19'd7,19'd1,-19'd44,-19'd12,19'd42,-19'd39,-19'd9,-19'd4,19'd15,19'd19,19'd8,19'd9,-19'd28,-19'd18,-19'd19,19'd49,-19'd25,19'd5,-19'd18,19'd3,19'd14,19'd3,19'd28,-19'd17,19'd14,-19'd40,19'd37,-19'd1,19'd1,19'd49,19'd39,19'd14,-19'd35,-19'd21,-19'd27,19'd37,19'd35,19'd33,-19'd25,-19'd48,-19'd10,-19'd40,19'd25,19'd18,19'd43,19'd48,19'd0,-19'd44,-19'd22,19'd47,19'd47,19'd1,19'd14,19'd43,19'd23,-19'd17,-19'd3,19'd29,19'd39,19'd21,-19'd38,-19'd28,19'd13,-19'd16,-19'd37,-19'd22,19'd36,-19'd6,-19'd15,-19'd10,19'd0,-19'd40,-19'd13,-19'd36,-19'd29,19'd47,19'd44,-19'd47,-19'd6,19'd19,19'd46,-19'd41,19'd20,-19'd27,19'd14,19'd9,19'd36,19'd25,-19'd42,19'd47,19'd15,19'd47,-19'd28,19'd49,19'd46,19'd15,19'd14,19'd15,19'd37,-19'd20,-19'd1,19'd47,-19'd32,-19'd11,-19'd8,-19'd7,-19'd13,19'd37,19'd11,-19'd22,-19'd10,-19'd46,-19'd40,19'd11,19'd25,19'd9,-19'd19,-19'd18,-19'd41,-19'd42,19'd21,-19'd22,-19'd33,-19'd30,19'd27,-19'd28,19'd23,19'd44,19'd49,19'd1,19'd23,19'd4,19'd36,19'd37,-19'd31,-19'd19,-19'd34,19'd28,19'd21,19'd28,19'd16,-19'd11,-19'd4,19'd40,19'd10,-19'd1,19'd9,-19'd27,19'd44,-19'd24,-19'd31,19'd35,19'd8,19'd32,-19'd49,-19'd13,-19'd6,-19'd39,19'd37,19'd42,19'd19,19'd30,-19'd37,-19'd6,19'd41,-19'd17,19'd1,19'd47,-19'd48,19'd28,19'd49,19'd1,-19'd36,19'd2,-19'd2,-19'd11,-19'd33,-19'd43,19'd32,19'd29,-19'd9,19'd7,19'd37,-19'd8,19'd31,19'd15,19'd19,19'd10,-19'd42,19'd34,19'd12,19'd46,19'd44,19'd0,19'd5,19'd28,-19'd11,19'd6,19'd1,-19'd50,19'd45,-19'd42,-19'd3,19'd16,19'd45,-19'd12,-19'd27,-19'd38,-19'd13,-19'd47,-19'd24,-19'd27,19'd15,-19'd25,19'd46,19'd45,-19'd22,-19'd3,-19'd22,19'd49,19'd30,-19'd6,-19'd47,-19'd9,-19'd31,-19'd21,19'd45,-19'd5,19'd1,-19'd18,-19'd29,19'd1,-19'd23,19'd10,19'd37,-19'd26,19'd28,19'd15,-19'd4,19'd20,19'd21,-19'd20,-19'd44,19'd21,-19'd12,19'd10,19'd42,19'd32,19'd49,-19'd39,-19'd39,-19'd18,19'd6,-19'd21,-19'd39,19'd29,-19'd2,19'd48,19'd47,19'd38,-19'd41,-19'd37,-19'd2,-19'd24,-19'd43,-19'd7,-19'd3,-19'd23,-19'd18,19'd16,19'd50,19'd18,-19'd19,19'd21,19'd18,-19'd43,19'd9,-19'd49,19'd14,-19'd40,-19'd18,19'd13,19'd2,-19'd25,19'd23,19'd48,19'd47,-19'd23,19'd5,19'd21,-19'd28,-19'd13,19'd4,19'd17,19'd5,-19'd6,19'd21,19'd43,-19'd12,-19'd48,19'd8,-19'd14,19'd0,-19'd22,19'd35,-19'd13,19'd12,19'd3,19'd2,-19'd17,19'd30,19'd39,19'd40,19'd46,19'd37,19'd34,-19'd48,19'd5,-19'd34,19'd24,19'd7,19'd10,-19'd31,-19'd33,19'd43,19'd21,19'd32,19'd50,-19'd25,19'd5,19'd46,19'd23,-19'd4,19'd1,-19'd28,-19'd29,19'd1,19'd7,19'd43,-19'd2,19'd22,-19'd50,-19'd44,19'd17,19'd25,-19'd11,19'd24,-19'd32,-19'd7,19'd49,19'd21,19'd28,-19'd49,-19'd18,-19'd9,-19'd44,-19'd5,-19'd31,-19'd37,-19'd38,-19'd34,-19'd47,-19'd18,-19'd25,19'd3,19'd45,19'd24,19'd44,-19'd4,19'd21,-19'd29,-19'd2,19'd47,-19'd25,-19'd48,19'd23,-19'd40,19'd31,-19'd33,19'd36,-19'd49,-19'd25,-19'd4,19'd4,19'd30,19'd43,-19'd47,19'd7,-19'd44,19'd11,-19'd1,-19'd47,-19'd39,19'd30,19'd31,-19'd50,19'd1,-19'd7,-19'd36,-19'd8,19'd47,-19'd34,19'd15,19'd43,-19'd29,19'd9,19'd47,19'd27,19'd12,19'd39,19'd22,19'd18,19'd18,19'd1,19'd22,19'd16,-19'd11,-19'd15,19'd30,-19'd29,-19'd7,19'd49,-19'd4,-19'd10,19'd45,-19'd8,19'd3,19'd49,19'd20,-19'd24,-19'd8,-19'd32,-19'd23,19'd0,-19'd18,-19'd36,-19'd34,-19'd13,19'd17,19'd44,-19'd12,19'd47,19'd13,-19'd35,-19'd10,19'd35,-19'd12,-19'd27,19'd26,-19'd31,-19'd43,19'd13,19'd11,-19'd16,19'd38,-19'd32,-19'd37,-19'd15,19'd1,-19'd46,19'd35,-19'd6,19'd45,-19'd19,19'd30,19'd1,19'd26,19'd6,-19'd46,-19'd21,19'd42,19'd36,-19'd32,-19'd37,-19'd38,19'd48,-19'd45,-19'd49,-19'd11,19'd39,-19'd20,-19'd39,19'd43,-19'd49,-19'd11,-19'd38,-19'd30,-19'd28,-19'd33,-19'd41,19'd36,19'd25,19'd21,19'd33,19'd18,-19'd5,19'd43,-19'd31,-19'd25,19'd5,19'd7,19'd0,19'd11,19'd25,-19'd10,19'd1,19'd35,-19'd15,19'd43,19'd1,19'd0,19'd39,19'd15,19'd21,19'd10,-19'd11,19'd45,-19'd44,-19'd35,19'd42,19'd39,19'd3,19'd45,-19'd25,19'd49,-19'd48,19'd9,-19'd32,-19'd32,19'd43,-19'd34,-19'd6,19'd44,-19'd40,-19'd4,-19'd12,-19'd43,19'd31,19'd10,-19'd31,19'd23,19'd14,19'd47,19'd35,19'd45,-19'd49,19'd25,-19'd40,19'd3,-19'd7,-19'd35,-19'd39,19'd41,19'd10,-19'd50,-19'd7,19'd29,19'd36,-19'd32,19'd10,19'd15,-19'd43,19'd30,-19'd28,19'd46,19'd26,-19'd40,19'd5,-19'd1,19'd6,-19'd19,-19'd18,-19'd39,19'd16,19'd29,-19'd18,-19'd29,-19'd21,-19'd49,-19'd28,-19'd16,19'd33,19'd21,-19'd47,-19'd10,19'd15,19'd26,19'd5,-19'd28,19'd0,19'd41,-19'd50,-19'd37,19'd32,19'd41,19'd13,-19'd8,19'd0,19'd1,19'd10,-19'd3,19'd2,19'd35,19'd45,19'd50,-19'd16,-19'd37,19'd20,-19'd3,-19'd7,19'd35,-19'd19,19'd45,19'd45,19'd47,19'd20,19'd41,-19'd35,19'd25,19'd2,19'd37,-19'd38,19'd10,19'd46,-19'd18,19'd37,19'd43,19'd13,-19'd31,-19'd9,-19'd16,19'd4,-19'd33,19'd16,-19'd44,-19'd43,-19'd22,19'd11,-19'd4,-19'd30,19'd35,-19'd23
		};
		
	end
	



endmodule