module Top(opcode, out);
input [2:0]opcode;
output [7:0]out;

////YOUR CODE/////////

endmodule