module Top(a, b, c, d);
input [1:0] a,b,c;
output [2:0]d;

///Your code////

endmodule
