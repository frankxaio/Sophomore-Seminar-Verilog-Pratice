module Top(sel,out);

input [1:0]sel;
output [3:0]out;

////YOUR CODE/////////

endmodule