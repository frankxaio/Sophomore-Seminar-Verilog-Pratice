module matrix_mutiply2(input [5999:0] image,
                       input [5999:0] weight,
                       input [299:0] Bias,
                       output reg [2999:0] Result); // 30*10*10
    
    reg [29:0] A1 [0:9][0:19];
    reg [29:0] B1 [0:19][0:9];
    reg [29:0] Bias_reg [0:9];
    reg [29:0] Res1 [0:9][0:9];
    
    integer i,j,k;
    
    always@ (image or weight) begin
        //We convert the 1D arrays into 2D
        {
        A1[0][0],A1[0][1],A1[0][2],A1[0][3],A1[0][4],A1[0][5],A1[0][6],A1[0][7],A1[0][8],A1[0][9],A1[0][10],A1[0][11],A1[0][12],A1[0][13],A1[0][14],A1[0][15],A1[0][16],A1[0][17],A1[0][18],A1[0][19],A1[1][0],A1[1][1],A1[1][2],A1[1][3],A1[1][4],A1[1][5],A1[1][6],A1[1][7],A1[1][8],A1[1][9],A1[1][10],A1[1][11],A1[1][12],A1[1][13],A1[1][14],A1[1][15],A1[1][16],A1[1][17],A1[1][18],A1[1][19],A1[2][0],A1[2][1],A1[2][2],A1[2][3],A1[2][4],A1[2][5],A1[2][6],A1[2][7],A1[2][8],A1[2][9],A1[2][10],A1[2][11],A1[2][12],A1[2][13],A1[2][14],A1[2][15],A1[2][16],A1[2][17],A1[2][18],A1[2][19],A1[3][0],A1[3][1],A1[3][2],A1[3][3],A1[3][4],A1[3][5],A1[3][6],A1[3][7],A1[3][8],A1[3][9],A1[3][10],A1[3][11],A1[3][12],A1[3][13],A1[3][14],A1[3][15],A1[3][16],A1[3][17],A1[3][18],A1[3][19],A1[4][0],A1[4][1],A1[4][2],A1[4][3],A1[4][4],A1[4][5],A1[4][6],A1[4][7],A1[4][8],A1[4][9],A1[4][10],A1[4][11],A1[4][12],A1[4][13],A1[4][14],A1[4][15],A1[4][16],A1[4][17],A1[4][18],A1[4][19],A1[5][0],A1[5][1],A1[5][2],A1[5][3],A1[5][4],A1[5][5],A1[5][6],A1[5][7],A1[5][8],A1[5][9],A1[5][10],A1[5][11],A1[5][12],A1[5][13],A1[5][14],A1[5][15],A1[5][16],A1[5][17],A1[5][18],A1[5][19],A1[6][0],A1[6][1],A1[6][2],A1[6][3],A1[6][4],A1[6][5],A1[6][6],A1[6][7],A1[6][8],A1[6][9],A1[6][10],A1[6][11],A1[6][12],A1[6][13],A1[6][14],A1[6][15],A1[6][16],A1[6][17],A1[6][18],A1[6][19],A1[7][0],A1[7][1],A1[7][2],A1[7][3],A1[7][4],A1[7][5],A1[7][6],A1[7][7],A1[7][8],A1[7][9],A1[7][10],A1[7][11],A1[7][12],A1[7][13],A1[7][14],A1[7][15],A1[7][16],A1[7][17],A1[7][18],A1[7][19],A1[8][0],A1[8][1],A1[8][2],A1[8][3],A1[8][4],A1[8][5],A1[8][6],A1[8][7],A1[8][8],A1[8][9],A1[8][10],A1[8][11],A1[8][12],A1[8][13],A1[8][14],A1[8][15],A1[8][16],A1[8][17],A1[8][18],A1[8][19],A1[9][0],A1[9][1],A1[9][2],A1[9][3],A1[9][4],A1[9][5],A1[9][6],A1[9][7],A1[9][8],A1[9][9],A1[9][10],A1[9][11],A1[9][12],A1[9][13],A1[9][14],A1[9][15],A1[9][16],A1[9][17],A1[9][18],A1[9][19]
        } = image;
        {
        B1[0][0],B1[0][1],B1[0][2],B1[0][3],B1[0][4],B1[0][5],B1[0][6],B1[0][7],B1[0][8],B1[0][9],B1[1][0],B1[1][1],B1[1][2],B1[1][3],B1[1][4],B1[1][5],B1[1][6],B1[1][7],B1[1][8],B1[1][9],B1[2][0],B1[2][1],B1[2][2],B1[2][3],B1[2][4],B1[2][5],B1[2][6],B1[2][7],B1[2][8],B1[2][9],B1[3][0],B1[3][1],B1[3][2],B1[3][3],B1[3][4],B1[3][5],B1[3][6],B1[3][7],B1[3][8],B1[3][9],B1[4][0],B1[4][1],B1[4][2],B1[4][3],B1[4][4],B1[4][5],B1[4][6],B1[4][7],B1[4][8],B1[4][9],B1[5][0],B1[5][1],B1[5][2],B1[5][3],B1[5][4],B1[5][5],B1[5][6],B1[5][7],B1[5][8],B1[5][9],B1[6][0],B1[6][1],B1[6][2],B1[6][3],B1[6][4],B1[6][5],B1[6][6],B1[6][7],B1[6][8],B1[6][9],B1[7][0],B1[7][1],B1[7][2],B1[7][3],B1[7][4],B1[7][5],B1[7][6],B1[7][7],B1[7][8],B1[7][9],B1[8][0],B1[8][1],B1[8][2],B1[8][3],B1[8][4],B1[8][5],B1[8][6],B1[8][7],B1[8][8],B1[8][9],B1[9][0],B1[9][1],B1[9][2],B1[9][3],B1[9][4],B1[9][5],B1[9][6],B1[9][7],B1[9][8],B1[9][9],B1[10][0],B1[10][1],B1[10][2],B1[10][3],B1[10][4],B1[10][5],B1[10][6],B1[10][7],B1[10][8],B1[10][9],B1[11][0],B1[11][1],B1[11][2],B1[11][3],B1[11][4],B1[11][5],B1[11][6],B1[11][7],B1[11][8],B1[11][9],B1[12][0],B1[12][1],B1[12][2],B1[12][3],B1[12][4],B1[12][5],B1[12][6],B1[12][7],B1[12][8],B1[12][9],B1[13][0],B1[13][1],B1[13][2],B1[13][3],B1[13][4],B1[13][5],B1[13][6],B1[13][7],B1[13][8],B1[13][9],B1[14][0],B1[14][1],B1[14][2],B1[14][3],B1[14][4],B1[14][5],B1[14][6],B1[14][7],B1[14][8],B1[14][9],B1[15][0],B1[15][1],B1[15][2],B1[15][3],B1[15][4],B1[15][5],B1[15][6],B1[15][7],B1[15][8],B1[15][9],B1[16][0],B1[16][1],B1[16][2],B1[16][3],B1[16][4],B1[16][5],B1[16][6],B1[16][7],B1[16][8],B1[16][9],B1[17][0],B1[17][1],B1[17][2],B1[17][3],B1[17][4],B1[17][5],B1[17][6],B1[17][7],B1[17][8],B1[17][9],B1[18][0],B1[18][1],B1[18][2],B1[18][3],B1[18][4],B1[18][5],B1[18][6],B1[18][7],B1[18][8],B1[18][9],B1[19][0],B1[19][1],B1[19][2],B1[19][3],B1[19][4],B1[19][5],B1[19][6],B1[19][7],B1[19][8],B1[19][9]
        } = weight;
        {
        Bias_reg[0] ,Bias_reg[1] ,Bias_reg[2] ,Bias_reg[3] ,Bias_reg[4] ,Bias_reg[5] ,Bias_reg[6] ,Bias_reg[7] ,Bias_reg[8] ,Bias_reg[9]
        } = Bias;
        {
        Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[0][4],Res1[0][5],Res1[0][6],Res1[0][7],Res1[0][8],Res1[0][9],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[1][4],Res1[1][5],Res1[1][6],Res1[1][7],Res1[1][8],Res1[1][9],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[2][4],Res1[2][5],Res1[2][6],Res1[2][7],Res1[2][8],Res1[2][9],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3],Res1[3][4],Res1[3][5],Res1[3][6],Res1[3][7],Res1[3][8],Res1[3][9],Res1[4][0],Res1[4][1],Res1[4][2],Res1[4][3],Res1[4][4],Res1[4][5],Res1[4][6],Res1[4][7],Res1[4][8],Res1[4][9],Res1[5][0],Res1[5][1],Res1[5][2],Res1[5][3],Res1[5][4],Res1[5][5],Res1[5][6],Res1[5][7],Res1[5][8],Res1[5][9],Res1[6][0],Res1[6][1],Res1[6][2],Res1[6][3],Res1[6][4],Res1[6][5],Res1[6][6],Res1[6][7],Res1[6][8],Res1[6][9],Res1[7][0],Res1[7][1],Res1[7][2],Res1[7][3],Res1[7][4],Res1[7][5],Res1[7][6],Res1[7][7],Res1[7][8],Res1[7][9],Res1[8][0],Res1[8][1],Res1[8][2],Res1[8][3],Res1[8][4],Res1[8][5],Res1[8][6],Res1[8][7],Res1[8][8],Res1[8][9],Res1[9][0],Res1[9][1],Res1[9][2],Res1[9][3],Res1[9][4],Res1[9][5],Res1[9][6],Res1[9][7],Res1[9][8],Res1[9][9]
        } = 3000'd0;
        
        i = 0; j = 0; k = 0;
        
        for(i = 0;i<10;i = i+1) begin
            for(j = 0;j<10;j = j+1) begin
                for(k = 0;k<20;k = k+1) begin
                    Res1[i][j] = Res1[i][j]+ (A1[i][k]*B1[k][j]);
                end
                if (Res1[i][j][29] == 1)
                    Res1[i][j] = 0;
                else
                    Res1[i][j] = Res1[i][j] + Bias_reg[j];
            end
        end
        // Turn 2D array into 1D
        Result = {
        Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[0][4],Res1[0][5],Res1[0][6],Res1[0][7],Res1[0][8],Res1[0][9],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[1][4],Res1[1][5],Res1[1][6],Res1[1][7],Res1[1][8],Res1[1][9],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[2][4],Res1[2][5],Res1[2][6],Res1[2][7],Res1[2][8],Res1[2][9],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3],Res1[3][4],Res1[3][5],Res1[3][6],Res1[3][7],Res1[3][8],Res1[3][9],Res1[4][0],Res1[4][1],Res1[4][2],Res1[4][3],Res1[4][4],Res1[4][5],Res1[4][6],Res1[4][7],Res1[4][8],Res1[4][9],Res1[5][0],Res1[5][1],Res1[5][2],Res1[5][3],Res1[5][4],Res1[5][5],Res1[5][6],Res1[5][7],Res1[5][8],Res1[5][9],Res1[6][0],Res1[6][1],Res1[6][2],Res1[6][3],Res1[6][4],Res1[6][5],Res1[6][6],Res1[6][7],Res1[6][8],Res1[6][9],Res1[7][0],Res1[7][1],Res1[7][2],Res1[7][3],Res1[7][4],Res1[7][5],Res1[7][6],Res1[7][7],Res1[7][8],Res1[7][9],Res1[8][0],Res1[8][1],Res1[8][2],Res1[8][3],Res1[8][4],Res1[8][5],Res1[8][6],Res1[8][7],Res1[8][8],Res1[8][9],Res1[9][0],Res1[9][1],Res1[9][2],Res1[9][3],Res1[9][4],Res1[9][5],Res1[9][6],Res1[9][7],Res1[9][8],Res1[9][9]
        };
    end
    
endmodule
