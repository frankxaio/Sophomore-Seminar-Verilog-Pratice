module Top (
	input [9:0] image [49:0]

);

always @( *) begin
	for (

    
end