module Top(a, b, sum,cout);
input [2:0]a,b;
output [2:0]sum,cout;

////YOUR CODE/////////

endmodule