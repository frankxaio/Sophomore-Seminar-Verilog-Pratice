module Top(clk,rst,plus,sub,out,seg7);

input	clk,rst,plus,sub;
output	[3:0]out;
output	[7:0] seg7;

////YOUR CODE/////////

endmodule