module Top(a, b, out);
input [3:0]a,b;
output [4:0]out;

////YOUR CODE/////////

endmodule