module Top(rst,clk,out,seg7);

input	clk,rst;
output	[3:0]out;
output	[7:0] seg7;

////YOUR CODE/////////

endmodule