module Maxmin (
    // input signals
    in_num,
    in_valid,
    rst_n,
    clk,

    // output signals
    out_valid,
    out_max,
    out_min
);

  //---------------------------------------------------------------------
  //   INPUT AND OUTPUT DECLARATION                         
  //---------------------------------------------------------------------


  //---------------------------------------------------------------------
  //   LOGIC DECLARATION
  //---------------------------------------------------------------------


  //---------------------------------------------------------------------
  //   Your design                        
  //---------------------------------------------------------------------



endmodule
