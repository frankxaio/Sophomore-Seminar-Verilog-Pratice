module Top(rst, clk, a, b, out, seg7);
input clk,rst;
input [3:0]a,b;
output [1:0]out;
output [7:0]seg7;

////YOUR CODE/////////

endmodule